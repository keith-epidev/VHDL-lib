function char2int(arg : character) return natural is
	begin
	return character'pos(arg);
end char2int;
